'
.include lib/bc847blp.mod

vcc 1 0  DC  3
Q1 1 2 3 bc847blp
Q2 2 1 3 bc847blp
L1 1 2 1u
C1 1 2 100p
R1 3 0 1K
C2 2 4 1n
R2 4 0 3K

.width out=140
.option rstray
.plot tran v 4 v 2
.tran 1n 300n

