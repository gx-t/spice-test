'
.include lib/bc847blp.mod
.include lib/bc857blp.mod

V1 1 0  DC 5

Q1 2 3 4 bc847blp
Q2 5 2 1 bc857blp
Q3 5 8 0 bc847blp
Q4 8 3 4 bc857blp

R1 5 0 10K
R2 4 5 100K
C2 4 7 1u
R5 7 0 10K

R3 1 3 51K
R4 3 0 51K
V2 6 0 AC 1
C1 6 3 1u


.width out=140
.option rstray

.print op v 4 v 5
.op


.print ac v 6 v 5
.ac 10 100e3 1e3
