'
.include 'lib/irl2505.spi'

V1 1 0 dc 5

XQ1 3 2 0 irl2505
R1 1 3 0.1

V2 4 0 pulse 0 5 10u 0 0 10u 300u
R2 4 2 300


.width out=140
.option rstray

.print tran v 4 i R1 i R2 v 2

.tran 1u 30u

