'
* Impedance

V2(1 0) sin (freq=100e6 ampl=1) AC 1
Rs(1 2) 50

C1(2, 0) 30p
L1(2, 3) 82nH
C2(3, 0) 30p

Rl(3, 0) 50

.width out=120
.option rstray

.print ac vdb(3) z(3)
.ac 88Meg 250Meg 1Meg
