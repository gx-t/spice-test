'
.include lib/LM741.MOD

V1 1 0 15V
V2 2 0 -15V
XOP 3 4 1 2 4 LM741/NS
V3 3 0 AC 4.5

.width out=140
.option rstray

.print op v 4 v 1 v 2
.op

.print ac vdb 4
.ac 100K 3Meg * 1.01

.plot ac v 4
.ac 100K 3Meg * 1.1

