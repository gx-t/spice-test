'
.include lib/bc847blp.mod

V1 vcc 0 DC  3
Q1 out base 0 bc847blp
R1 out base 1Meg
R2 out vcc 4.7k

C1 base rc 1000p
C2 out rc 1000p
R3 rc in 100K
V2 in 0 AC 1

.print op v out
.op

.width out=140
.option rstray

.print ac vdb out
.ac 200 2100 * 1.01

.plot ac vdb out
.ac 200 2100 * 1.01

