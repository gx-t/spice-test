'
.include lib/2sc3356.mod
.include lib/ss9018g.mod
.include lib/BFR520.MOD

* FM transmitter output amplifier

V1(vcc 0) DC 5

V2(1, 0) sin (freq=101.5Meg ampl=14m) AC 14m

R1(1,in) 50
C1(in,q1_b) 330p

Q1(q1_c,q1_b,0) BFR520
R1(q1_c,q1_b) 47K
L1(q1_c,vcc) 80n
C2(q1_c,out) 47p
C3(out,0) 68p
Rout(out,0) 50

.width out=120
.option rstray

.print op i(q1)
.op

.print ac z(q1_b) z(out) v(out) p(Rout) v(q1_c)
.ac 88Meg 108Meg 1Meg

.plot tran v(out)(-1,1)
.tran 1u 4u 0.2n

'.plot fourier v(7)
'.fourier 88Meg 1G 1Meg

