'
.include 'lib/irl2505.spi'

V1 1 0 dc 5

XQ1 3 2 0 irl2505
R1 1 3 0.1

V2 4 0 PULSE 0 10 1n 1n 1n 500n 1000n
R2 4 2 1


.width out=140
.option rstray

.print tran i R1 i R2 v 2

.tran 20n 1000n

