'
.include 'lib/irl2505.spi'

V1 1 0 dc 5

XQ1 3 2 0 irl2505
R1 1 3 0.1

'TC4420 2.5ohm, 25ns, 25ns
V2 4 0 pulse 0 5 10u 25n 25n 10u 300u
R2 4 2 2.5


.width out=140
.option rstray

.print tran v 4 i R1 i R2 v 2

.tran 10u 10.2u 5n
.tran 20u 20.2u 5n

.plot tran i R1

.tran 10u 10.2u 5n
.tran 20u 20.2u 5n

